module control #(
	parameter RESET_ADDR = 32'h00000000
)(
	input wire [5:0] opcode,
	input wire [2:0] funct3,
	input wire [6:0] funct7,
	output wire [1:0] alu_op,
	output wire 

);




endmodule