module execute #(
	parameter RESET_ADDR = 32'h00000000
);

// Most of this instantiates our ALU we already made





endmodule