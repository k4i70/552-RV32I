module hart #(
    // After reset, the program counter (PC) should be initialized to this
    // address and start executing instructions from there.
    parameter RESET_ADDR = 32'h00000000
) (
    // Global clock.
    input  wire        i_clk,
    // Synchronous active-high reset.
    input  wire        i_rst,
    // Instruction fetch goes through a read only instruction memory (imem)
    // port. The port accepts a 32-bit address (e.g. from the program counter)
    // per cycle and combinationally returns a 32-bit instruction word. This
    // is not representative of a realistic memory interface; it has been
    // modeled as more similar to a DFF or SRAM to simplify phase 3. In
    // later phases, you will replace this with a more realistic memory.
    //
    // 32-bit read address for the instruction memory. This is expected to be
    // 4 byte aligned - that is, the two LSBs should be zero.
    output wire [31:0] o_imem_raddr,
    // Instruction word fetched from memory, available on the same cycle.
    input  wire [31:0] i_imem_rdata,
    // Data memory accesses go through a separate read/write data memory (dmem)
    // that is shared between read (load) and write (stored). The port accepts
    // a 32-bit address, read or write enable, and mask (explained below) each
    // cycle. Reads are combinational - values are available immediately after
    // updating the address and asserting read enable. Writes occur on (and
    // are visible at) the next clock edge.
    //
    // Read/write address for the data memory. This should be 32-bit aligned
    // (i.e. the two LSB should be zero). See `o_dmem_mask` for how to perform
    // half-word and byte accesses at unaligned addresses.
    output wire [31:0] o_dmem_addr,
    // When asserted, the memory will perform a read at the aligned address
    // specified by `i_addr` and return the 32-bit word at that address
    // immediately (i.e. combinationally). It is illegal to assert this and
    // `o_dmem_wen` on the same cycle.
    output wire        o_dmem_ren,
    // When asserted, the memory will perform a write to the aligned address
    // `o_dmem_addr`. When asserted, the memory will write the bytes in
    // `o_dmem_wdata` (specified by the mask) to memory at the specified
    // address on the next rising clock edge. It is illegal to assert this and
    // `o_dmem_ren` on the same cycle.
    output wire        o_dmem_wen,
    // The 32-bit word to write to memory when `o_dmem_wen` is asserted. When
    // write enable is asserted, the byte lanes specified by the mask will be
    // written to the memory word at the aligned address at the next rising
    // clock edge. The other byte lanes of the word will be unaffected.
    output wire [31:0] o_dmem_wdata,
    // The dmem interface expects word (32 bit) aligned addresses. However,
    // WISC-25 supports byte and half-word loads and stores at unaligned and
    // 16-bit aligned addresses, respectively. To support this, the access
    // mask specifies which bytes within the 32-bit word are actually read
    // from or written to memory.
    //
    // To perform a half-word read at address 0x00001002, align `o_dmem_addr`
    // to 0x00001000, assert `o_dmem_ren`, and set the mask to 0b1100 to
    // indicate that only the upper two bytes should be read. Only the upper
    // two bytes of `i_dmem_rdata` can be assumed to have valid data; to
    // calculate the final value of the `lh[u]` instruction, shift the rdata
    // word right by 16 bits and sign/zero extend as appropriate.
    //
    // To perform a byte write at address 0x00002003, align `o_dmem_addr` to
    // `0x00002000`, assert `o_dmem_wen`, and set the mask to 0b1000 to
    // indicate that only the upper byte should be written. On the next clock
    // cycle, the upper byte of `o_dmem_wdata` will be written to memory, with
    // the other three bytes of the aligned word unaffected. Remember to shift
    // the value of the `sb` instruction left by 24 bits to place it in the
    // appropriate byte lane.
    output wire [ 3:0] o_dmem_mask,
    // The 32-bit word read from data memory. When `o_dmem_ren` is asserted,
    // this will immediately reflect the contents of memory at the specified
    // address, for the bytes enabled by the mask. When read enable is not
    // asserted, or for bytes not set in the mask, the value is undefined.
    input  wire [31:0] i_dmem_rdata,
	// The output `retire` interface is used to signal to the testbench that
    // the CPU has completed and retired an instruction. A single cycle
    // implementation will assert this every cycle; however, a pipelined
    // implementation that needs to stall (due to internal hazards or waiting
    // on memory accesses) will not assert the signal on cycles where the
    // instruction in the writeback stage is not retiring.
    //
    // Asserted when an instruction is being retired this cycle. If this is
    // not asserted, the other retire signals are ignored and may be left invalid.
    output wire        o_retire_valid,
    // The 32 bit instruction word of the instrution being retired. This
    // should be the unmodified instruction word fetched from instruction
    // memory.
    output wire [31:0] o_retire_inst,
    // Asserted if the instruction produced a trap, due to an illegal
    // instruction, unaligned data memory access, or unaligned instruction
    // address on a taken branch or jump.
    output wire        o_retire_trap,
    // Asserted if the instruction is an `ebreak` instruction used to halt the
    // processor. This is used for debugging and testing purposes to end
    // a program.
    output wire        o_retire_halt,
    // The first register address read by the instruction being retired. If
    // the instruction does not read from a register (like `lui`), this
    // should be 5'd0.
    output wire [ 4:0] o_retire_rs1_raddr,
    // The second register address read by the instruction being retired. If
    // the instruction does not read from a second register (like `addi`), this
    // should be 5'd0.
    output wire [ 4:0] o_retire_rs2_raddr,
    // The first source register data read from the register file (in the
    // decode stage) for the instruction being retired. If rs1 is 5'd0, this
    // should also be 32'd0.
    output wire [31:0] o_retire_rs1_rdata,
    // The second source register data read from the register file (in the
    // decode stage) for the instruction being retired. If rs2 is 5'd0, this
    // should also be 32'd0.
    output wire [31:0] o_retire_rs2_rdata,
    // The destination register address written by the instruction being
    // retired. If the instruction does not write to a register (like `sw`),
    // this should be 5'd0.
    output wire [ 4:0] o_retire_rd_waddr,
    // The destination register data written to the register file in the
    // writeback stage by this instruction. If rd is 5'd0, this field is
    // ignored and can be treated as a don't care.
    output wire [31:0] o_retire_rd_wdata,
    // The current program counter of the instruction being retired - i.e.
    // the instruction memory address that the instruction was fetched from.
    output wire [31:0] o_retire_pc,
    // the next program counter after the instruction is retired. For most
    // instructions, this is `o_retire_pc + 4`, but must be the branch or jump
    // target for *taken* branches and jumps.
    output wire [31:0] o_retire_next_pc

`ifdef RISCV_FORMAL
    ,`RVFI_OUTPUTS,
`endif
);
    // Fill in your implementation here.

    // Intermediate signals
    wire [6:0] opcode;
    wire [31:0] address_in;
    wire [2:0] funct3;
    wire [2:0] mem_funct3;
    wire [6:0] funct7;
    wire [3:0] branch_op;
    wire [31:0] o_rs1_data;
    wire [31:0] o_rs2_data;
    wire [4:0] rd;
    wire [31:0] o_immediate;
    wire [5:0] o_format;
    wire [2:0] alu_op;
    wire [1:0] reg_write_source_op;
    wire [31:0] rs1_data;
    wire [31:0] rs2_data;
    wire [31:0] immediate;
    wire [31:0] alu_result;
    wire [31:0] branch_out;
    wire [31:0] WriteData;
    wire [4:0] rd_out;
    wire [31:0] mem_raddr;
    wire [4:0] rs1_raddr;
    wire [4:0] rs2_raddr;
    wire [3:0] dmem_mask_base;
    wire [31:0] load_data;

    wire mem_write, reg_write, alu_src_op, pc_src_op, o_eq, o_slt, i_sub, i_unsigned, i_arith;
    wire reg_write_wb, jalr_op, alu_pc_op, mem_read;

    // Gate register writes with valid to prevent writes during the reset cycle
    wire reg_write_wb_safe = reg_write_wb & o_retire_valid;

    assign mem_funct3 = i_imem_rdata[14:12];

    


    // Split into pipelined stages 
    // Have specific files for each stage. 
    // Piece of advice from people who have taken the class before, split into a bunch of small subfiles
    // So most of the code is probably just connecting all the subfiles


    /** Instruction Fetch **/
    fetch i_fetch (
        .i_clk(i_clk),
        .i_rst(i_rst),
        .address_in(address_in), 
        .o_mem_raddr(o_imem_raddr),
        .o_retire_valid(o_retire_valid)
    );



    /** Instruction Decode **/
    decode i_decode (
        .i_clk(i_clk),
        .i_rst(i_rst),
        .i_instr(i_imem_rdata),
        .opcode(opcode),
        .rd(rd),
        .o_immediate(immediate),
        .o_format(o_format),
        .alu_op(alu_op),
        .branch_op(branch_op),
        .mem_write(mem_write),
        .reg_write_source_op(reg_write_source_op),
        .reg_write(reg_write),
        .alu_src_op(alu_src_op),
        .pc_src_op(pc_src_op),
        .o_dmem_mask(dmem_mask_base),
        .i_sub(i_sub),
        .i_unsigned(i_unsigned),
        .i_arith(i_arith),
        .o_rs1_rdata(rs1_data),
        .o_rs2_rdata(rs2_data),
        .reg_write_wb(reg_write_wb_safe),
        .i_rd_waddr(rd_out),
        .i_rd_wdata(WriteData),
        .rs1_raddr(rs1_raddr),
        .rs2_raddr(rs2_raddr),
        .jalr_op(jalr_op),
        .alu_pc_op(alu_pc_op),
        .mem_read(mem_read)
    );
        

    /** Execute **/
    execute i_execute (
        .pc_src_op(pc_src_op),
        .alu_src_op(alu_src_op),
        .alu_op(alu_op),
        .rs1_data(rs1_data),
        .rs2_data(rs2_data),
        .immediate(immediate),
        .alu_result(alu_result),
        .o_eq(o_eq),
        .o_slt(o_slt),
        .i_sub(i_sub),
        .i_unsigned(i_unsigned),
        .i_arith(i_arith),
        .branch_op(branch_op),
        .branch_out(branch_out),
        .jalr_op(jalr_op),
        .alu_pc_op(alu_pc_op),
        .PC(o_imem_raddr)
    );



    /** Memory Access **/
    memoryAccess i_memoryAccess (
        .mem_write(mem_write),
        .alu_result(alu_result), 
        .rs2_data(rs2_data),
        .o_dmem_addr(o_dmem_addr), 
        .o_dmem_wdata(o_dmem_wdata),
        .o_dmem_ren(o_dmem_ren),
        .o_dmem_wen(o_dmem_wen),
        .i_dmem_rdata(i_dmem_rdata),
        .o_dmem_mask(o_dmem_mask),
        .dmem_mask_base(dmem_mask_base),
        .mem_read(mem_read),
        .funct3(mem_funct3),
        .i_unsigned(i_unsigned),
        .o_load_data(load_data)
    );


    /** Writeback **/
    writeback i_writeback (
        .RegWrite(reg_write),
        .rd(rd),
        .PC(o_imem_raddr),
        .branch_out(branch_out),
        .ALUResult(alu_result),
        .ReadData(load_data),
        .MemtoReg(reg_write_source_op),
        .pc_src_op(pc_src_op),
        .rd_out(rd_out),
        .WriteData(WriteData),
        .reg_write_wb(reg_write_wb),
        .current_PC(address_in),
        .jalr_op(jalr_op)
    );


    // Declare retire signals and connect with assigns
    assign o_retire_inst = i_imem_rdata;
    assign o_retire_trap = 1'b0; 
    assign o_retire_halt = (i_imem_rdata == 32'h00100073); // Ebreak instruction
    assign o_retire_rs1_raddr = i_imem_rdata[19:15];
    assign o_retire_rs2_raddr = i_imem_rdata[24:20];
    assign o_retire_rs1_rdata = rs1_data;
    assign o_retire_rs2_rdata = rs2_data;
    assign o_retire_rd_waddr = rd_out;
    assign o_retire_rd_wdata = WriteData;
    assign o_retire_pc = o_imem_raddr;
    assign o_retire_next_pc = address_in;


endmodule

`default_nettype wire
