module execute #(
	parameter RESET_ADDR = 32'h00000000
);





endmodule